`define clock_sensor_data_width              8
`define window_sensor_data_width             8
`define daylight_sensor_data_width           8
`define motion_sensor_data_width             8
`define security_sensor_data_width           8
`define temperature_sensor_data_width        8
`define ac_cool_data_width                   8
`define heating_system_on_off_data_width     8
`define door_motion_sensor_data_width        4
`define light_threshold                      128
`define temp_threshold                       128
